module fifo #(
    //parameters
)(
    //io
);

    // stuffz
endmodule

