module uart #(
  //params
  
)(
  //io
    
);
  
endmodule

